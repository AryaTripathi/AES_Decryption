module Inverse_sbox(s_in, s_out);
    
input  [7:0] s_in;
output reg [7:0] s_out; 
always @(*)
begin
case (s_in)	

 8'h00 : s_out =  8'h16;
 8'h01 : s_out =  8'hbb;
 8'h02 : s_out =  8'h54;
 8'h03 : s_out =  8'hb0;
 8'h04 : s_out =  8'h0f;
 8'h05 : s_out =  8'h2d;
 8'h06 : s_out =  8'h99;
 8'h07 : s_out =  8'h41;
 8'h08 : s_out =  8'h68;
 8'h09 : s_out =  8'h42;
 8'h0A : s_out =  8'he6;
 8'h0B : s_out =  8'hbf;
 8'h0C : s_out =  8'h0d;
 8'h0D : s_out =  8'h89;
 8'h0E : s_out =  8'ha1;
 8'h0F : s_out =  8'h8c;
 8'h10 : s_out =  8'hdf;
 8'h11 : s_out =  8'h28;
 8'h12 : s_out =  8'h55;
 8'h13 : s_out =  8'hce;
 8'h14 : s_out =  8'he9;
 8'h15 : s_out =  8'h87;
 8'h16 : s_out =  8'h1e;
 8'h17 : s_out =  8'h9b;
 8'h18 : s_out =  8'h94;
 8'h19 : s_out =  8'h8e;
 8'h1A : s_out =  8'hd9;
 8'h1B : s_out =  8'h69;
 8'h1C : s_out =  8'h11;
 8'h1D : s_out =  8'h98;
 8'h1E : s_out =  8'hf8;
 8'h1F : s_out =  8'he1;
 8'h20 : s_out =  8'h9e;
 8'h21 : s_out =  8'h1d;
 8'h22 : s_out =  8'hc1;
 8'h23 : s_out =  8'h86;
 8'h24 : s_out =  8'hb9;
 8'h25 : s_out =  8'h57;
 8'h26 : s_out =  8'h35;
 8'h27 : s_out =  8'h61;
 8'h28 : s_out =  8'h0e;
 8'h29 : s_out =  8'hf6;
 8'h2A : s_out =  8'h03;
 8'h2B : s_out =  8'h48;
 8'h2C : s_out =  8'h66;
 8'h2D : s_out =  8'hb5;
 8'h2E : s_out =  8'h3e;
 8'h2F : s_out =  8'h70;
 8'h30 : s_out =  8'h8a;
 8'h31 : s_out =  8'h8b;
 8'h32 : s_out =  8'hbd;
 8'h33 : s_out =  8'h4b;
 8'h34 : s_out =  8'h1f;
 8'h35 : s_out =  8'h74;
 8'h36 : s_out =  8'hdd;
 8'h37 : s_out =  8'he8;
 8'h38 : s_out =  8'hc6;
 8'h39 : s_out =  8'hb4;
 8'h3A : s_out =  8'ha6;
 8'h3B : s_out =  8'h1c;
 8'h3C : s_out =  8'h2e;
 8'h3D : s_out =  8'h25;
 8'h3E : s_out =  8'h78;
 8'h3F : s_out =  8'hba;
 8'h40 : s_out =  8'h08;
 8'h41 : s_out =  8'hae;
 8'h42 : s_out =  8'h7a;
 8'h43 : s_out =  8'h65;
 8'h44 : s_out =  8'hea;
 8'h45 : s_out =  8'hf4;
 8'h46 : s_out =  8'h56;
 8'h47 : s_out =  8'h6c;
 8'h48 : s_out =  8'ha9;
 8'h49 : s_out =  8'h4e;
 8'h4A : s_out =  8'hd5;
 8'h4B : s_out =  8'h8d;
 8'h4C : s_out =  8'h6d;
 8'h4D : s_out =  8'h37;
 8'h4E : s_out =  8'hc8;
 8'h4F : s_out =  8'he7;
 8'h50 : s_out =  8'h79;
 8'h51 : s_out =  8'he4;
 8'h52 : s_out =  8'h95;
 8'h53 : s_out =  8'h91;
 8'h54 : s_out =  8'h62;
 8'h55 : s_out =  8'hac;
 8'h56 : s_out =  8'hd3;
 8'h57 : s_out =  8'hc2;
 8'h58 : s_out =  8'h5c;
 8'h59 : s_out =  8'h24;
 8'h5A : s_out =  8'h06;
 8'h5B : s_out =  8'h49;
 8'h5C : s_out =  8'h0a;
 8'h5D : s_out =  8'h3a;
 8'h5E : s_out =  8'h32;
 8'h5F : s_out =  8'he0;
 8'h60 : s_out =  8'hdb;
 8'h61 : s_out =  8'h0b;
 8'h62 : s_out =  8'h5e;
 8'h63 : s_out =  8'hde;
 8'h64 : s_out =  8'h14;
 8'h65 : s_out =  8'hb8;
 8'h66 : s_out =  8'hee;
 8'h67 : s_out =  8'h46;
 8'h68 : s_out =  8'h88;
 8'h69 : s_out =  8'h90;
 8'h6A : s_out =  8'h2a;
 8'h6B : s_out =  8'h22;
 8'h6C : s_out =  8'hdc;
 8'h6D : s_out =  8'h4f;
 8'h6E : s_out =  8'h81;
 8'h6F : s_out =  8'h60;
 8'h70 : s_out =  8'h73;
 8'h71 : s_out =  8'h19;
 8'h72 : s_out =  8'h5d;
 8'h73 : s_out =  8'h64;
 8'h74 : s_out =  8'h3d;
 8'h75 : s_out =  8'h7e;
 8'h76 : s_out =  8'ha7;
 8'h77 : s_out =  8'hc4;
 8'h78 : s_out =  8'h17;
 8'h79 : s_out =  8'h44;
 8'h7A : s_out =  8'h97;
 8'h7B : s_out =  8'h5f;
 8'h7C : s_out =  8'hec;
 8'h7D : s_out =  8'h13;
 8'h7E : s_out =  8'h0c;
 8'h7F : s_out =  8'hcd;
 8'h80 : s_out =  8'hd2;
 8'h81 : s_out =  8'hf3;
 8'h82 : s_out =  8'hff;
 8'h83 : s_out =  8'h10;
 8'h84 : s_out =  8'h21;
 8'h85 : s_out =  8'hda;
 8'h86 : s_out =  8'hb6;
 8'h87 : s_out =  8'hbc;
 8'h88 : s_out =  8'hf5;
 8'h89 : s_out =  8'h38;
 8'h8A : s_out =  8'h9d;
 8'h8B : s_out =  8'h92;
 8'h8C : s_out =  8'h8f;
 8'h8D : s_out =  8'h40;
 8'h8E : s_out =  8'ha3;
 8'h8F : s_out =  8'h51;
 8'h90 : s_out =  8'ha8;
 8'h91 : s_out =  8'h9f;
 8'h92 : s_out =  8'h3c;
 8'h93 : s_out =  8'h50;
 8'h94 : s_out =  8'h7f;
 8'h95 : s_out =  8'h02;
 8'h96 : s_out =  8'hf9;
 8'h97 : s_out =  8'h45;
 8'h98 : s_out =  8'h85;
 8'h99 : s_out =  8'h33;
 8'h9A : s_out =  8'h4d;
 8'h9B : s_out =  8'h43;
 8'h9C : s_out =  8'hfb;
 8'h9D : s_out =  8'haa;
 8'h9E : s_out =  8'hef;
 8'h9F : s_out =  8'hd0;
 8'hA0 : s_out =  8'hcf;
 8'hA1 : s_out =  8'h58;
 8'hA2 : s_out =  8'h4c;
 8'hA3 : s_out =  8'h4a;
 8'hA4 : s_out =  8'h39;
 8'hA5 : s_out =  8'hbe;
 8'hA6 : s_out =  8'hcb;
 8'hA7 : s_out =  8'h6a;
 8'hA8 : s_out =  8'h5b;
 8'hA9 : s_out =  8'hb1;
 8'hAA : s_out =  8'hfc;
 8'hAB : s_out =  8'h20;
 8'hAC : s_out =  8'hed;
 8'hAD : s_out =  8'h00;
 8'hAE : s_out =  8'hd1;
 8'hAF : s_out =  8'h53;
 8'hB0 : s_out =  8'h84;
 8'hB1 : s_out =  8'h2f;
 8'hB2 : s_out =  8'he3;
 8'hB3 : s_out =  8'h29;
 8'hB4 : s_out =  8'hb3;
 8'hB5 : s_out =  8'hd6;
 8'hB6 : s_out =  8'h3b;
 8'hB7 : s_out =  8'h52;
 8'hB8 : s_out =  8'ha0;
 8'hB9 : s_out =  8'h5a;
 8'hBA : s_out =  8'h6e;
 8'hBB : s_out =  8'h1b;
 8'hBC : s_out =  8'h1a;
 8'hBD : s_out =  8'h2c;
 8'hBE : s_out =  8'h83;
 8'hBF : s_out =  8'h09;
 8'hC0 : s_out =  8'h75;
 8'hC1 : s_out =  8'hb2;
 8'hC2 : s_out =  8'h27;
 8'hC3 : s_out =  8'heb;
 8'hC4 : s_out =  8'he2;
 8'hC5 : s_out =  8'h80;
 8'hC6 : s_out =  8'h12;
 8'hC7 : s_out =  8'h07;
 8'hC8 : s_out =  8'h9a;
 8'hC9 : s_out =  8'h05;
 8'hCA : s_out =  8'h96;
 8'hCB : s_out =  8'h18;
 8'hCC : s_out =  8'hc3;
 8'hCD : s_out =  8'h23;
 8'hCE : s_out =  8'hc7;
 8'hCF : s_out =  8'h04;
 8'hD0 : s_out =  8'h15;
 8'hD1 : s_out =  8'h31;
 8'hD2 : s_out =  8'hd8;
 8'hD3 : s_out =  8'h71;
 8'hD4 : s_out =  8'hf1;
 8'hD5 : s_out =  8'he5;
 8'hD6 : s_out =  8'ha5;
 8'hD7 : s_out =  8'h34;
 8'hD8 : s_out =  8'hcc;
 8'hD9 : s_out =  8'hf7;
 8'hDA : s_out =  8'h3f;
 8'hDB : s_out =  8'h36;
 8'hDC : s_out =  8'h26;
 8'hDD : s_out =  8'h93;
 8'hDE : s_out =  8'hfd;
 8'hDF : s_out =  8'hb7;
 8'hE0 : s_out =  8'hc0;
 8'hE1 : s_out =  8'h72;
 8'hE2 : s_out =  8'ha4;
 8'hE3 : s_out =  8'h9c;
 8'hE4 : s_out =  8'haf;
 8'hE5 : s_out =  8'ha2;
 8'hE6 : s_out =  8'hd4;
 8'hE7 : s_out =  8'had;
 8'hE8 : s_out =  8'hf0;
 8'hE9 : s_out =  8'h47;
 8'hEA : s_out =  8'h59;
 8'hEB : s_out =  8'hfa;
 8'hEC : s_out =  8'h7d;
 8'hED : s_out =  8'hc9;
 8'hEE : s_out =  8'h82;
 8'hEF : s_out =  8'hca;
 8'hF0 : s_out =  8'h76;
 8'hF1 : s_out =  8'hab;
 8'hF2 : s_out =  8'hd7;
 8'hF3 : s_out =  8'hfe;
 8'hF4 : s_out =  8'h2b;
 8'hF5 : s_out =  8'h67;
 8'hF6 : s_out =  8'h01;
 8'hF7 : s_out =  8'h30;
 8'hF8 : s_out =  8'hc5;
 8'hF9 : s_out =  8'h6f;
 8'hFA : s_out =  8'h6b;
 8'hFB : s_out =  8'hf2;
 8'hFC : s_out =  8'h7b;
 8'hFD : s_out =  8'h77;
 8'hFE : s_out =  8'h7c;
 8'hFF : s_out =  8'h63;
 
endcase
end
endmodule
